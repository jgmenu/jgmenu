Terminal,^term(bash)
Filhanterare,pcmanfm
Webbläsare,firefox
Textredigerare,^term(vim)
^sep()
Tillbehör,^checkout(accessories)
^sep()
Platser,^pipe(jgmenu_run places)
^sep()
Hjälp och Information,^checkout(help)
^sep()
Lås skärmen,i3lock-fancy -p

^tag(accessories)
Post,:
Meddelande,:
Fildelning,:
Skärmbild,:

^tag(help)
Hjälp,:
Information,:
